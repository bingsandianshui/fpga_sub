library verilog;
use verilog.vl_types.all;
entity LTC1744_T01_tb is
end LTC1744_T01_tb;
