module find_start();

endmodule
